op3 <= op1 and op2;
