op2 <= (31 downto 30 => op1(31)) & op1(31 downto 2);