op3 <= std_logic_vector(signed(op1) + signed(op2));
op4 <= std_logic_vector(signed(op1) - signed(op2));
