-- megafunction wizard: %ROM: 1-PORT%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: altsyncram 

-- ============================================================
-- File Name: crc_tta_stratix_altera_onchip_rom_comp.vhd
-- Megafunction Name(s):
--          altsyncram
--
-- Simulation Library Files(s):
--          
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 8.0 Build 215 05/29/2008 SJ Full Version
-- ************************************************************


--Copyright (C) 1991-2008 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


library ieee;
use ieee.std_logic_1164.all;

library altera_mf;
use altera_mf.all;

entity ENTITY_STR_altera_onchip_rom_comp is
  generic (
    init_file_g  : string  := "init_data.mif";
    dev_family_g : string  := "Cyclone II";
    addrw_g      : integer := 10;
    dataw_g      : integer := 32);
  port (
    address : in  std_logic_vector (addrw_g-1 downto 0);
    clken   : in  std_logic;
    clock   : in  std_logic;
    q       : out std_logic_vector (dataw_g-1 downto 0));
end ENTITY_STR_altera_onchip_rom_comp;


architecture SYN of ENTITY_STR_altera_onchip_rom_comp is

  signal sub_wire0 : std_logic_vector (dataw_g-1 downto 0);

  component altsyncram
    generic (
      clock_enable_input_a   : string;
      clock_enable_output_a  : string;
      init_file              : string;
      intended_device_family : string;
      lpm_hint               : string;
      lpm_type               : string;
      numwords_a             : natural;
      operation_mode         : string;
      outdata_aclr_a         : string;
      outdata_reg_a          : string;
      widthad_a              : natural;
      width_a                : natural;
      width_byteena_a        : natural
      );
    port (
      clocken0  : in  std_logic;
      clock0    : in  std_logic;
      address_a : in  std_logic_vector (addrw_g-1 downto 0);
      q_a       : out std_logic_vector (dataw_g-1 downto 0)
      );
  end component;

begin
  q <= sub_wire0(dataw_g-1 downto 0);

  altsyncram_component : altsyncram
    generic map (
      clock_enable_input_a   => "NORMAL",
      clock_enable_output_a  => "BYPASS",
      init_file              => init_file_g,
      intended_device_family => dev_family_g,
      lpm_hint               => "ENABLE_RUNTIME_MOD=NO",
      lpm_type               => "altsyncram",
      numwords_a             => 2**addrw_g,
      operation_mode         => "ROM",
      outdata_aclr_a         => "NONE",
      outdata_reg_a          => "UNREGISTERED",
      widthad_a              => addrw_g,
      width_a                => dataw_g,
      width_byteena_a        => 1
      )
    port map (
      clocken0  => clken,
      clock0    => clock,
      address_a => address,
      q_a       => sub_wire0
      );

end SYN;
