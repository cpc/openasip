load_data_32b <= rdata_out_1;
op2 <= load_data_32b;
