op2 <= op1(27 downto 0) & "0000";