op3 <= std_logic_vector(unsigned(op1) rem unsigned(op2));