if op1 /= op2 then
  op3 <= '1';
else
  op3 <= '0';
end if;
