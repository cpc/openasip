op2 <= "0000" & op1(31 downto 4);