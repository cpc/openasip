op2 <= (31 downto 24 => op1(31)) & op1(31 downto 8);