op2 <= not op1(15) & op1(14 downto 0);
