-- Copyright (c) 2002-2012 Tampere University.
--
-- This file is part of TTA-Based Codesign Environment (TCE).
-- 
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the "Software"),
-- to deal in the Software without restriction, including without limitation
-- the rights to use, copy, modify, merge, publish, distribute, sublicense,
-- and/or sell copies of the Software, and to permit persons to whom the
-- Software is furnished to do so, subject to the following conditions:
-- 
-- The above copyright notice and this permission notice shall be included in
-- all copies or substantial portions of the Software.
-- 
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
-- IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
-- FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
-- AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
-- LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING
-- FROM, OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER
-- DEALINGS IN THE SOFTWARE.
---------------------------------------------------------------------------------
-- Title      : Register File for TTA
-- Project    : FlexDSP
-------------------------------------------------------------------------------
-- Original arch:
-- VHDL Architecture RF_lib.rf_4wr_4rd_always_1.symbol
--
-- Created:  10:55:33 11/22/05
--          by - tpitkane.tpitkane (elros)
--          at - 10:55:33 11/22/05
--
-- Generated by Mentor Graphics' HDL Designer(TM) 2004.1 (Build 41)
---------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author   Description
-- 8.6.2012    1.0      eskoo    Created
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
library work;
use work.util.all;

entity rf_4wr_7rd_always_1 is
  generic(
    dataw   : integer := 32;
    rf_size : integer := 4
    );
  port(
    clk      : in  std_logic;
    rstx     : in std_logic;    
    glock    : in  std_logic;
    -- read ports
    r1load   : in  std_logic;
    r1opcode : in  std_logic_vector(bit_width(rf_size)-1 downto 0);
    r1data   : out std_logic_vector(dataw-1 downto 0);
    r2load   : in  std_logic;
    r2opcode : in  std_logic_vector(bit_width(rf_size)-1 downto 0);
    r2data   : out std_logic_vector(dataw-1 downto 0);
    r3load   : in  std_logic;
    r3opcode : in  std_logic_vector(bit_width(rf_size)-1 downto 0);
    r3data   : out std_logic_vector(dataw-1 downto 0);
    r4load   : in  std_logic;
    r4opcode : in  std_logic_vector(bit_width(rf_size)-1 downto 0);
    r4data   : out std_logic_vector(dataw-1 downto 0);
    r5load   : in  std_logic;
    r5opcode : in  std_logic_vector(bit_width(rf_size)-1 downto 0);
    r5data   : out std_logic_vector(dataw-1 downto 0);
    r6load   : in  std_logic;
    r6opcode : in  std_logic_vector(bit_width(rf_size)-1 downto 0);
    r6data   : out std_logic_vector(dataw-1 downto 0);
    r7load   : in  std_logic;
    r7opcode : in  std_logic_vector(bit_width(rf_size)-1 downto 0);
    r7data   : out std_logic_vector(dataw-1 downto 0);
    -- writer ports
    t1data   : in std_logic_vector(dataw-1 downto 0);
    t1load   : in std_logic;
    t1opcode : in std_logic_vector(bit_width(rf_size)-1 downto 0);
    t2data   : in std_logic_vector(dataw-1 downto 0);
    t2load   : in std_logic;
    t2opcode : in std_logic_vector(bit_width(rf_size)-1 downto 0);
    t3data   : in std_logic_vector(dataw-1 downto 0);
    t3load   : in std_logic;
    t3opcode : in std_logic_vector(bit_width(rf_size)-1 downto 0);
    t4data   : in std_logic_vector(dataw-1 downto 0);
    t4load   : in std_logic;
    t4opcode : in std_logic_vector(bit_width(rf_size)-1 downto 0)
    );

-- Declarations

end rf_4wr_7rd_always_1;
---------------------------------------------------------------------------------
-- Title      : Register File for TTA
-- Project    : FlexDSP
-------------------------------------------------------------------------------
--Original arch:
-- VHDL Architecture RF_lib.rf_4wr_4rd_always_1.rtl
--
-- Created:  10:55:33 11/22/05
--          by - tpitkane.tpitkane (elros)
--          at - 10:55:33 11/22/05
--
-- Generated by Mentor Graphics' HDL Designer(TM) 2004.1 (Build 41)
---------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author   Description
-- 8.6.2012    1.0    eskoo    Created
---------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
library work;
use work.util.all;
architecture rtl of rf_4wr_7rd_always_1 is

  -- Architecture declarations
  type    reg_type is array (natural range <>) of std_logic_vector(dataw-1 downto 0);
  subtype rf_index is integer range 0 to rf_size-1;
  signal  reg : reg_type (rf_size-1 downto 0);

begin

  -----------------------------------------------------------------
  Input : process (clk, rstx)
    -----------------------------------------------------------------

    -- Process declarations
    variable opc : integer;


  begin
    -- Asynchronous Reset
    if (rstx = '0') then
      -- Reset Actions
      for idx in (reg'length-1) downto 0 loop
        reg(idx) <= (others => '0');
      end loop;  -- idx

    elsif (clk'event and clk = '1') then
      if glock = '0' then
        if t1load = '1' then
          opc      := conv_integer(unsigned(t1opcode));
          reg(opc) <= t1data;
        end if;
        if t2load = '1' then
          opc      := conv_integer(unsigned(t2opcode));
          reg(opc) <= t2data;
        end if;
        if t3load = '1' then
          opc      := conv_integer(unsigned(t3opcode));
          reg(opc) <= t3data;
        end if;
        if t4load = '1' then
          opc      := conv_integer(unsigned(t4opcode));
          reg(opc) <= t4data;
        end if;
      end if;
    end if;
  end process Input;

  -----------------------------------------------------------------
  --output : PROCESS (glock, r1load, r1opcode, r2load, r2opcode, r3load, r3opcode, r4load, r4opcode, reg, rstx)
  -----------------------------------------------------------------

  r1data <= reg(conv_integer(unsigned(r1opcode)));
  r2data <= reg(conv_integer(unsigned(r2opcode)));
  r3data <= reg(conv_integer(unsigned(r3opcode)));
  r4data <= reg(conv_integer(unsigned(r4opcode)));
  r5data <= reg(conv_integer(unsigned(r5opcode)));
  r6data <= reg(conv_integer(unsigned(r6opcode)));
  r7data <= reg(conv_integer(unsigned(r7opcode)));
  
end rtl;
