op2 <= op1(29 downto 0) & "00";