op2 <= op1(15 downto 0) & X"0000";