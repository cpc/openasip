op3 <= op1 or op2;
