op4 <= std_logic_vector(resize(unsigned(op1) + unsigned(op2) * unsigned(op3), op4'length));
