op3 <= std_logic_vector(resize(unsigned(op1) * unsigned(op2), op3'length));
