op3 <= std_logic_vector(shift_right(signed(op1), to_integer(unsigned(op2(4 downto 0)))));
