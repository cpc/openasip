op2 <= "0" & op1(31 downto 1);