op2 <= '0' & op1(14 downto 0);
