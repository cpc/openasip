op3 <= std_logic_vector(rotate_right(unsigned(op1), to_integer(signed(op2))));
