op2 <= "00" & op1(31 downto 2);