op3 <= op1 xor op2;
