if unsigned(op1) > unsigned(op2) then
  op3 <= op1;
else
  op3 <= op2;
end if;
