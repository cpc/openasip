if op3(0) = '1' then
    op4 <= op1;
else
    op4 <= op2;
end if;