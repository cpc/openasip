op2 <= std_logic_vector(resize(signed(op1), 32));
