avalid_in_1 <= '1';
aaddr_in_1 <= op1(addrw_c-1 downto 0);
awren_in_1 <= '0';
