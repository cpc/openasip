avalid_in_1 <= '1';
awren_in_1 <= '1';
aaddr_in_1 <= op1(addrw_c-1 downto 0);
adata_in_1 <= op2;
astrb_in_1 <= "1111";
