op3 <= std_logic_vector(signed(op1) + signed(op2));
