if signed(op1) < signed(op2) then
  op3 <= '0';
else
  op3 <= '1';
end if;
