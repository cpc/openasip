if unsigned(op1) < unsigned(op2) then
  op3 <= '0';
else
  op3 <= '1';
end if;
