op3 <= std_logic_vector(resize(shift_right(resize(signed(op1), 33) * signed(resize(unsigned(op2), 33)), 32), 32));