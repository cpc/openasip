op2 <= op1(31) & op1(31 downto 1);