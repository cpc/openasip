if signed(op1) < signed(op2) then
  op3 <= '1';
else
  op3 <= '0';
end if;
