op3 <= std_logic_vector(rotate_left(unsigned(op1), to_integer(unsigned(op2))));
