---------------------------------------------------------------------------------
-- Title        : File for TTA
-- Project    : FlexDSP
-------------------------------------------------------------------------------
--
-- VHDL Architecture RF_lib.rf_1wr_1rd_always_1.symbol
--
-- Created:  10:55:31 11/22/05
--          by - tpitkane.tpitkane (elros)
--          at - 10:55:31 11/22/05
--
-- Generated by Mentor Graphics' HDL Designer(TM) 2004.1 (Build 41)
---------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author   Description
-- 11/22/05      1.0     tpitkane   Created
-------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;
USE work.util.all;

ENTITY rf_1wr_0rd_always_1 IS
   GENERIC( 
      dataw   : integer := 32;
      rf_size : integer := 8
   );
   PORT( 
      clk      : IN     std_logic;
      glock    : IN     std_logic;
      rstx     : IN     std_logic;
      t1data   : IN     std_logic_vector (dataw-1 DOWNTO 0);
      t1load   : IN     std_logic;
      t1opcode : IN     std_logic_vector ( bit_width(rf_size)-1 DOWNTO 0 );
      guard    : out    std_logic_vector ( rf_size-1 DOWNTO 0)
   );

-- Declarations

END rf_1wr_0rd_always_1 ;
---------------------------------------------------------------------------------
-- Title        : File for TTA
-- Project    : FlexDSP
-------------------------------------------------------------------------------
--
-- VHDL Architecture RF_lib.rf_1wr_1rd_always_1.rtl
--
-- Created:  10:55:31 11/22/05
--          by - tpitkane.tpitkane (elros)
--          at - 10:55:31 11/22/05
--
-- Generated by Mentor Graphics' HDL Designer(TM) 2004.1 (Build 41)
---------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author   Description
-- 11/22/05      1.0     tpitkane   Created
---------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;
ARCHITECTURE rtl OF rf_1wr_0rd_always_1 IS

   -- Architecture declarations
   type   reg_type is array (natural range <>) of std_logic_vector(dataw-1 downto 0 );
   subtype rf_index is integer range 0 to rf_size-1;
   signal reg    : reg_type (rf_size-1 downto 0);

   signal t1data_orred : std_logic_vector(0 downto 0);
BEGIN

   -----------------------------------------------------------------
   input : PROCESS (clk, rstx)
   -----------------------------------------------------------------

   -- Process declarations
   variable opc : integer;


   BEGIN
      -- Asynchronous Reset
      IF (rstx = '0') THEN
         -- Reset Actions
         for idx in (reg'length-1) downto 0 loop
           reg(idx) <= (others => '0');
         end loop;  -- idx

      ELSIF (clk'EVENT AND clk = '1') THEN
         IF glock = '0' THEN
            IF t1load = '1' THEN
               opc := conv_integer(unsigned(t1opcode));
               reg(opc) <= t1data;
            END IF;
         END IF;
      END IF;
   END PROCESS input;

   OR_t1data: process (t1data)
     variable orred_t1data : std_logic_vector(0 downto 0);
   begin  -- process OR_t1data
     orred_t1data := "0";
     for i in t1data'range loop
       orred_t1data := t1data(i downto i) or (orred_t1data);
     end loop;
     t1data_orred <= orred_t1data;
       
   end process OR_t1data;

     
   guard_process: process (t1load,t1opcode,t1data_orred,rstx)
     variable opc : integer;
     
   begin  -- process guard
     if rstx = '0' then
       guard <= (others => '0');
     else
       if glock = '0' then
         if t1load = '1' then
           opc := conv_integer(unsigned(t1opcode));
           guard(opc downto opc) <= t1data_orred; 
         end if;
       end if;
     end if;
     
   end process guard_process;
END rtl;
