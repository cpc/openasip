op2 <= X"0000" & op1(31 downto 16);