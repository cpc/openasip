op2 <= X"00" & op1(31 downto 8);