op3 <= std_logic_vector(resize(shift_right(unsigned(op1) * unsigned(op2), 32), 32));