op2 <= debug_lock_count_in(32-1 downto 0);