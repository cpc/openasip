if unsigned(op1) > unsigned(op2) then
  op3 <= '1';
else
  op3 <= '0';
end if;
