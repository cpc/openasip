-- AXI4-Lite master
m_axi_awaddr   => m_axi_awaddr,
m_axi_awvalid  => m_axi_awvalid,
m_axi_awready  => m_axi_awready,
m_axi_awprot   => m_axi_awprot,
m_axi_wvalid   => m_axi_wvalid,
m_axi_wready   => m_axi_wready,
m_axi_wdata    => m_axi_wdata,
m_axi_wstrb    => m_axi_wstrb,
m_axi_bvalid   => m_axi_bvalid,
m_axi_bready   => m_axi_bready,
m_axi_arvalid  => m_axi_arvalid,
m_axi_arready  => m_axi_arready,
m_axi_araddr   => m_axi_araddr,
m_axi_arprot   => m_axi_arprot,
m_axi_rdata    => m_axi_rdata,
m_axi_rvalid   => m_axi_rvalid,
m_axi_rready   => m_axi_rready,
