if signed(op1) > signed(op2) then
  op3 <= op2;
else
  op3 <= op1;
end if;
