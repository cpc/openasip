op2 <= op1(23 downto 0) & X"00";