op2 <= op1(30 downto 0) & "0";