op2 <= (31 downto 28 => op1(31)) & op1(31 downto 4);